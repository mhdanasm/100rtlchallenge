module B( input x,y, output z);
  xnor a1(z,x,y);
  
endmodule
